//------------------------------------------------------------------------------------------------------
// Company:        Xilinx & HES//SO hepia
// Engineer:       Xavier Paillard
// 
// Create Date:    08:49:58 01/29/2013 
// Design Name:    DVI
// Module Name:    PB_DVI_INIT
// Project Name:   DVI
// Target Devices: Xilinx SP605 - XC6SLX45T-3fpgg484
// Tool versions:  Xilinx ISE 14.3 - Windows 7 64bits
// Description:    This is a module for storing a program for the KCPSM3 (aka Pico-Blaze)
//                 The code is assembled as "pbt3" (should be pbt3 for spartan 3)
// Dependencies:   No
// Revision:       05-11-2004 Initial creation
//                 30-01-2013 File modified by Xavier Paillard, add simplification
//------------------------------------------------------------------------------------------------------

module PB_DVI_INIT
	(
	 CLK,        // Clock @ 125 MHz
	 ADDRESS,    // Read address
	 INSTRUCTION // Instruction bus
  );

	input	 CLK;
	input	 [9:0]  ADDRESS;
	output [17:0] INSTRUCTION;
	  
	RAMB16_S18_S18 rom
		(	
		 // Port A: Read Port
		 .CLKA(CLK),                 
		 .ADDRA(ADDRESS),            
		 .DIA(16'h0000),             
		 .DIPA(2'b00), 
		 .WEA(1'b0),
		 .DOA(INSTRUCTION[15:0]), 
		 .DOPA(INSTRUCTION[17:16]),
		 .ENA(1'b1), 
		 .SSRA(1'b0),
		 // port B: Load (write) port
		 .CLKB(1'b0), 
		 .ADDRB(10'b0000000000), 
		 .DIB(16'h0000), 
		 .DIPB(2'b00), 
		 .WEB(1'b0),
		 .DOB(), 
		 .DOPB(),
		 .ENB(1'b0), 
		 .SSRB(1'b0)
	  );	  

	// Init ROM with program
	defparam rom.INIT_00  = 256'h00740600054900740608052300740643051D007406090521E00200EC4001003E;
	defparam rom.INIT_01  = 256'h0104000A007406C0054901040032007406600536007406160534007406080533;
	defparam rom.INIT_02  = 256'h0074067005350074060805330074060C05330074061805480074061005480D14;
	defparam rom.INIT_03  = 256'hE00200ECA0005421CD015435CC01543DA80400AC00A1E003004DE00100010C14;
	defparam rom.INIT_04  = 256'h053400740606053300740600054900740608052300740643051D007406090521;
	defparam rom.INIT_05  = 256'h0074061005480D140104000A007406C0054901040032007406A0053600740626;
	defparam rom.INIT_06  = 256'hCC015473A80400AC00A1E003004DE00100010C14007406700535007406180548;
	defparam rom.INIT_07  = 256'h00B51860B400290100B085011850B400290100B0680200DCA000545DCD01546B;
	defparam rom.INIT_08  = 256'h00B51860B40000B01870B400290100B085011850B400290100B0680200DCA000;
	defparam rom.INIT_09  = 256'h00B06804B0004001600100B06803B00040006001B400290100B0680200DCA000;
	defparam rom.INIT_0A  = 256'h40ED00B808FF090140B808FF0900A00000B0C801680200DCB40029010091A000;
	defparam rom.INIT_0B  = 256'h000C00FA0A05C000000000010806010840ED00B8090140EDB000290100B80901;
	defparam rom.INIT_0C  = 256'hC000C002A001109054B9C10100FA0A05C0000008D800A001400000FA0A0AC000;
	defparam rom.INIT_0D  = 256'h00FA0A05C0000003A00000FA0A05C0000008490000FA0A0AC000000C00FA0A05;
	defparam rom.INIT_0E  = 256'h0A05C0000002A00000FA0A05C000000800FA0A05C000000200FA0A05C000000C;
	defparam rom.INIT_0F  = 256'hCB02CB0150FF2B01CB060B19A00000FA0A05C000000300FA0A05C000000C00FA;
	defparam rom.INIT_10  = 256'h8000A0005504C00100FA0AFA00FA0AFA00FA0AFA00FA0AFAA00054FACA0154FF;
	defparam rom.INIT_11  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_12  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_13  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_14  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_15  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_16  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_17  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_18  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_19  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_1F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_20  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_21  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_22  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_23  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_24  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_25  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_26  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_27  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_28  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_29  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_2F  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_30  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_31  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_32  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_33  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_34  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_35  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_36  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_37  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_38  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_39  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3A  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3B  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3C  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3D  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3E  = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INIT_3F  = 256'h410F000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INITP_00 = 256'hC9D273B773E20C30C0CC330C30C30C308B773E20C30C30C0CC330C30C30C308F;
	defparam rom.INITP_01 = 256'h5D4B232322C8C8C8C8B20C8C80DC80323288F39CF0C2C39EC93249CECB2749CE;
	defparam rom.INITP_02 = 256'h00000000000000000000000000000000000000000000000000000000EDCCCCB7;
	defparam rom.INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	defparam rom.INITP_07 = 256'hC000000000000000000000000000000000000000000000000000000000000000;

endmodule 