-- Top level for mandelbrot calculator
--  use : MandelbrotCounter, MandelbrotFSM & MandelbrotComplexCalculator

-- Progress:
--  - MandelbrotCounter           : [x] Compile, [ ] Test
--  - MandelbrotFSM               : [ ] Compile, [ ] Test
--  - MandelbrotComplexCalculator : [ ] Compile, [ ] Test
